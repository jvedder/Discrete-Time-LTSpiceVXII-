* Copyright (C) 2022 John Vedder. MIT License.
*
* Difference Block
.subckt diff out in1 in2
B1 out 0 V=v(in1) - v(in2)
.ends sum
